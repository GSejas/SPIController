`timescale 1ns / 1ps

module SPISegmentoControlado();


endmodule
